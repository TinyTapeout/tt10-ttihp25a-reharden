magic
tech sky130A
timestamp 1741564516
<< nwell >>
rect -66 149 720 320
rect -66 148 33 149
<< nmos >>
rect 109 27 142 98
rect 168 27 201 98
rect 384 27 404 70
rect 558 27 578 76
<< pmos >>
rect 109 167 142 243
rect 168 167 201 243
rect 384 200 404 243
rect 558 196 578 243
<< ndiff >>
rect 70 85 109 98
rect 70 38 80 85
rect 99 38 109 85
rect 70 27 109 38
rect 142 27 168 98
rect 201 79 243 98
rect 201 45 209 79
rect 228 45 243 79
rect 201 37 243 45
rect 273 62 384 70
rect 273 44 278 62
rect 295 44 384 62
rect 201 27 238 37
rect 273 27 384 44
rect 404 56 493 70
rect 404 38 471 56
rect 489 38 493 56
rect 404 27 493 38
rect 521 66 558 76
rect 521 33 531 66
rect 548 33 558 66
rect 521 27 558 33
rect 578 63 617 76
rect 578 44 591 63
rect 610 44 617 63
rect 578 27 617 44
<< pdiff >>
rect 70 242 109 243
rect 67 226 109 242
rect 67 179 77 226
rect 96 179 109 226
rect 67 168 109 179
rect 70 167 109 168
rect 142 167 168 243
rect 201 225 237 243
rect 273 225 384 243
rect 201 216 243 225
rect 201 182 210 216
rect 229 182 243 216
rect 273 207 277 225
rect 294 207 384 225
rect 273 200 384 207
rect 404 225 493 243
rect 404 207 472 225
rect 489 207 493 225
rect 404 200 493 207
rect 521 232 558 243
rect 521 202 531 232
rect 548 202 558 232
rect 201 174 243 182
rect 201 167 237 174
rect 521 196 558 202
rect 578 219 617 243
rect 578 201 589 219
rect 606 201 617 219
rect 578 196 617 201
<< ndiffc >>
rect 80 38 99 85
rect 209 45 228 79
rect 278 44 295 62
rect 471 38 489 56
rect 531 33 548 66
rect 591 44 610 63
<< pdiffc >>
rect 77 179 96 226
rect 210 182 229 216
rect 277 207 294 225
rect 472 207 489 225
rect 531 202 548 232
rect 589 201 606 219
<< poly >>
rect 109 243 142 256
rect 168 243 201 256
rect 384 243 404 256
rect 558 243 578 256
rect 109 149 142 167
rect 168 149 201 167
rect 109 142 145 149
rect 109 123 120 142
rect 138 123 145 142
rect 109 116 145 123
rect 168 142 205 149
rect 168 123 180 142
rect 198 123 205 142
rect 168 116 205 123
rect 384 119 404 200
rect 558 159 578 196
rect 499 152 585 159
rect 499 135 516 152
rect 533 135 585 152
rect 499 126 585 135
rect 109 98 142 116
rect 168 98 201 116
rect 367 114 417 119
rect 367 89 378 114
rect 404 89 417 114
rect 367 80 417 89
rect 384 70 404 80
rect 558 76 578 126
rect 109 14 142 27
rect 168 14 201 27
rect 384 14 404 27
rect 558 14 578 27
<< polycont >>
rect 120 123 138 142
rect 180 123 198 142
rect 516 135 533 152
rect 378 89 404 114
<< locali >>
rect 67 236 106 242
rect 67 173 73 236
rect 100 173 106 236
rect 445 237 500 243
rect 270 225 309 233
rect 201 216 243 225
rect 201 182 210 216
rect 229 182 243 216
rect 270 207 277 225
rect 294 207 309 225
rect 270 199 309 207
rect 445 203 454 237
rect 485 225 500 237
rect 489 207 500 225
rect 485 203 500 207
rect 270 198 297 199
rect 201 174 243 182
rect 276 174 297 198
rect 445 196 500 203
rect 521 232 554 241
rect 521 202 530 232
rect 552 202 554 232
rect 521 192 554 202
rect 581 219 632 225
rect 581 201 589 219
rect 606 201 632 219
rect 581 183 632 201
rect 67 168 106 173
rect 225 167 297 174
rect 111 142 147 150
rect 111 123 120 142
rect 138 123 147 142
rect 111 115 147 123
rect 171 142 207 150
rect 171 123 180 142
rect 198 123 207 142
rect 171 115 207 123
rect 226 148 233 167
rect 250 148 297 167
rect 226 143 297 148
rect 226 98 243 143
rect 72 89 106 95
rect 72 33 75 89
rect 102 33 106 89
rect 202 79 243 98
rect 202 72 209 79
rect 201 45 209 72
rect 228 45 243 79
rect 280 74 297 143
rect 507 152 545 155
rect 507 151 516 152
rect 533 151 545 152
rect 507 133 513 151
rect 534 133 545 151
rect 507 130 545 133
rect 367 114 417 119
rect 367 89 378 114
rect 404 109 417 114
rect 589 117 632 183
rect 589 109 619 117
rect 404 91 619 109
rect 404 89 417 91
rect 367 80 417 89
rect 201 37 243 45
rect 269 62 308 74
rect 269 44 278 62
rect 295 44 308 62
rect 269 39 308 44
rect 451 62 500 74
rect 72 30 106 33
rect 73 29 106 30
rect 451 35 463 62
rect 487 56 500 62
rect 489 38 500 56
rect 487 35 500 38
rect 451 27 500 35
rect 523 66 556 73
rect 589 72 619 91
rect 523 33 528 66
rect 550 33 556 66
rect 581 63 619 72
rect 581 44 591 63
rect 610 44 619 63
rect 581 37 619 44
rect 523 29 556 33
<< viali >>
rect 73 226 100 236
rect 73 179 77 226
rect 77 179 96 226
rect 96 179 100 226
rect 73 173 100 179
rect 454 225 485 237
rect 454 207 472 225
rect 472 207 485 225
rect 454 203 485 207
rect 530 202 531 232
rect 531 202 548 232
rect 548 202 552 232
rect 233 148 250 167
rect 75 85 102 89
rect 75 38 80 85
rect 80 38 99 85
rect 99 38 102 85
rect 75 33 102 38
rect 513 135 516 151
rect 516 135 533 151
rect 533 135 534 151
rect 513 133 534 135
rect 463 56 487 62
rect 463 38 471 56
rect 471 38 487 56
rect 463 35 487 38
rect 528 33 531 66
rect 531 33 548 66
rect 548 33 550 66
<< metal1 >>
rect 0 244 669 297
rect 67 236 106 244
rect 67 173 73 236
rect 100 173 106 236
rect 210 237 669 244
rect 210 233 454 237
rect 445 203 454 233
rect 485 233 669 237
rect 485 203 500 233
rect 445 196 500 203
rect 521 232 558 233
rect 521 202 530 232
rect 552 202 558 232
rect 521 194 558 202
rect 67 168 106 173
rect 225 170 256 172
rect 225 167 545 170
rect 225 148 233 167
rect 250 151 545 167
rect 250 149 513 151
rect 250 148 256 149
rect 225 145 256 148
rect 501 133 513 149
rect 534 149 545 151
rect 534 133 544 149
rect 501 126 544 133
rect 72 89 106 95
rect 72 70 75 89
rect 71 41 75 70
rect 69 33 75 41
rect 102 70 106 89
rect 102 33 107 70
rect 457 62 496 70
rect 457 35 463 62
rect 487 35 496 62
rect 457 33 496 35
rect 521 66 557 70
rect 521 33 528 66
rect 550 33 557 66
rect 0 -11 668 33
rect 0 -12 162 -11
<< labels >>
flabel metal1 483 -11 658 27 0 FreeSans 120 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 103 -11 278 27 0 FreeSans 120 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 304 -11 479 27 0 FreeSans 120 180 0 0 VGND
port 1 nsew ground bidirectional
flabel viali 513 133 534 151 0 FreeSans 120 0 0 0 X
flabel metal1 304 243 479 287 0 FreeSans 120 180 0 0 VPWR
port 2 nsew power bidirectional
flabel locali 233 149 250 168 0 FreeSans 120 0 0 0 X
flabel locali 174 117 206 147 0 FreeSans 120 0 0 0 B
port 5 nsew signal input
flabel locali 113 117 145 147 0 FreeSans 120 0 0 0 A
port 4 nsew signal input
flabel metal1 103 244 133 287 0 FreeSans 120 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal1 483 243 658 287 0 FreeSans 120 0 0 0 VPWR
port 2 nsew power bidirectional
flabel locali 595 123 626 152 0 FreeSans 120 0 0 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 670 272
string LEFclass CORE
string LEFsite unithd
string LEFsource USER
<< end >>
