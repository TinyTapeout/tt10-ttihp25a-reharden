VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO celem
  CLASS CORE ;
  FOREIGN celem ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.700 BY 2.720 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.720 0.300 1.060 0.950 ;
        RECT 0.730 0.290 1.060 0.300 ;
        RECT 4.510 0.270 5.000 0.740 ;
        RECT 5.230 0.290 5.560 0.730 ;
      LAYER met1 ;
        RECT 0.720 0.700 1.060 0.950 ;
        RECT 0.710 0.410 1.070 0.700 ;
        RECT 0.690 0.330 1.070 0.410 ;
        RECT 4.570 0.330 4.960 0.700 ;
        RECT 5.210 0.330 5.570 0.700 ;
        RECT 0.000 -0.110 6.680 0.330 ;
        RECT 0.000 -0.120 1.620 -0.110 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.670 1.680 1.060 2.420 ;
        RECT 4.450 1.960 5.000 2.430 ;
        RECT 5.210 1.920 5.540 2.410 ;
      LAYER met1 ;
        RECT 0.000 2.440 6.690 2.970 ;
        RECT 0.670 1.680 1.060 2.440 ;
        RECT 2.100 2.330 6.690 2.440 ;
        RECT 4.450 1.960 5.000 2.330 ;
        RECT 5.210 1.940 5.580 2.330 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.172000 ;
    ANTENNADIFFAREA 0.374400 ;
    PORT
      LAYER li1 ;
        RECT 5.810 1.830 6.320 2.250 ;
        RECT 3.670 1.090 4.170 1.190 ;
        RECT 5.890 1.170 6.320 1.830 ;
        RECT 5.890 1.090 6.190 1.170 ;
        RECT 3.670 0.910 6.190 1.090 ;
        RECT 3.670 0.800 4.170 0.910 ;
        RECT 5.890 0.720 6.190 0.910 ;
        RECT 5.810 0.370 6.190 0.720 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.485100 ;
    PORT
      LAYER li1 ;
        RECT 1.110 1.150 1.470 1.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.485100 ;
    PORT
      LAYER li1 ;
        RECT 1.710 1.150 2.070 1.500 ;
    END
  END B
  OBS
      LAYER nwell ;
        RECT -0.660 1.490 7.200 3.200 ;
        RECT -0.660 1.480 0.330 1.490 ;
      LAYER li1 ;
        RECT 2.010 1.740 2.430 2.250 ;
        RECT 2.700 1.990 3.090 2.330 ;
        RECT 2.700 1.980 2.970 1.990 ;
        RECT 2.760 1.740 2.970 1.980 ;
        RECT 2.250 1.670 2.970 1.740 ;
        RECT 2.260 1.430 2.970 1.670 ;
        RECT 2.260 0.980 2.430 1.430 ;
        RECT 2.020 0.720 2.430 0.980 ;
        RECT 2.800 0.740 2.970 1.430 ;
        RECT 5.070 1.300 5.450 1.550 ;
        RECT 2.010 0.370 2.430 0.720 ;
        RECT 2.690 0.390 3.080 0.740 ;
      LAYER met1 ;
        RECT 2.250 1.700 2.560 1.720 ;
        RECT 2.250 1.490 5.450 1.700 ;
        RECT 2.250 1.450 2.560 1.490 ;
        RECT 5.010 1.260 5.440 1.490 ;
  END
END celem
END LIBRARY

