magic
tech sky130A
magscale 1 2
timestamp 1740304500
<< metal1 >>
rect 15540 43560 15660 43580
rect 15540 43480 15560 43560
rect 15640 43480 15660 43560
rect 15540 35300 15660 43480
rect 15540 35220 15560 35300
rect 15640 35220 15660 35300
rect 15540 35200 15660 35220
rect 9520 31400 9700 31420
rect 9520 31100 9540 31400
rect 9680 31100 9700 31400
rect 9520 30640 9700 31100
rect 12220 31400 12420 31420
rect 12220 31100 12240 31400
rect 12400 31100 12420 31400
rect 12220 30640 12420 31100
rect 14980 31400 15180 31420
rect 14980 31100 15000 31400
rect 15160 31100 15180 31400
rect 14980 30620 15180 31100
rect 17720 31400 17920 31420
rect 17720 31100 17740 31400
rect 17900 31100 17920 31400
rect 17720 30620 17920 31100
rect 20920 31260 21120 31280
rect 20920 31100 20940 31260
rect 21100 31100 21120 31260
rect 20920 31095 21120 31100
rect 11640 28780 11840 29020
rect 11640 28320 11660 28780
rect 11820 28320 11840 28780
rect 11640 28300 11840 28320
rect 14340 28780 14540 29020
rect 14340 28320 14360 28780
rect 14520 28320 14540 28780
rect 14340 28300 14540 28320
rect 16460 28780 16660 28800
rect 16460 28320 16480 28780
rect 16640 28320 16660 28780
rect 16460 28310 16660 28320
rect 17100 28780 17300 29020
rect 17100 28320 17120 28780
rect 17280 28320 17300 28780
rect 16460 24500 16771 28310
rect 17100 28300 17300 28320
rect 19840 28780 20040 29020
rect 19840 28320 19860 28780
rect 20020 28320 20040 28780
rect 19840 28300 20040 28320
rect 20797 27520 21120 31095
rect 20797 27516 20938 27520
rect 22960 25280 25060 25480
rect 22960 25020 23160 25280
rect 22640 24820 23160 25020
rect 24860 25000 25060 25280
rect 16460 24400 17180 24500
rect 16460 24180 17140 24400
rect 22640 24360 22860 24820
rect 13410 22240 13420 23380
rect 13540 22240 13550 23380
rect 15400 22920 16420 23140
rect 15400 22891 16359 22920
rect 15400 21800 15689 22891
rect 9300 21780 15689 21800
rect 9300 21620 9320 21780
rect 9680 21620 15689 21780
rect 9300 21600 15689 21620
rect 9663 21551 15689 21600
rect 15579 21547 15689 21551
rect 24860 20240 25060 22280
rect 16010 20060 16020 20220
rect 17940 20060 17950 20220
rect 21080 20040 25060 20240
<< via1 >>
rect 15560 43480 15640 43560
rect 15560 35220 15640 35300
rect 9540 31100 9680 31400
rect 12240 31100 12400 31400
rect 15000 31100 15160 31400
rect 17740 31100 17900 31400
rect 20940 31100 21100 31260
rect 11660 28320 11820 28780
rect 14360 28320 14520 28780
rect 16480 28320 16640 28780
rect 17120 28320 17280 28780
rect 19860 28320 20020 28780
rect 13420 22240 13540 23380
rect 9320 21620 9680 21780
rect 16020 20060 17940 20220
<< metal2 >>
rect 14540 43820 14660 43840
rect 14540 43740 14560 43820
rect 14640 43740 14660 43820
rect 14540 37000 14660 43740
rect 15540 43560 15780 43580
rect 15540 43480 15560 43560
rect 15640 43480 15680 43560
rect 15760 43480 15780 43560
rect 15540 43460 15780 43480
rect 28160 42720 28300 42740
rect 21040 42620 28180 42720
rect 28280 42620 28300 42720
rect 21040 42600 28300 42620
rect 21040 42200 21160 42600
rect 28720 42200 28860 42220
rect 18980 42080 21160 42200
rect 23040 42100 28740 42200
rect 28840 42100 28860 42200
rect 28720 42080 28860 42100
rect 14540 36920 14560 37000
rect 14640 36920 14660 37000
rect 14540 36900 14660 36920
rect 15540 35300 15660 35320
rect 15540 35220 15560 35300
rect 15640 35220 15660 35300
rect 15540 34980 15660 35220
rect 15540 34900 15560 34980
rect 15640 34900 15660 34980
rect 15540 34880 15660 34900
rect 9540 31400 9680 31410
rect 9540 31090 9680 31100
rect 12240 31400 12400 31410
rect 12240 31090 12400 31100
rect 15000 31400 15160 31410
rect 15000 31090 15160 31100
rect 17740 31400 17900 31410
rect 21040 31270 21100 31880
rect 17740 31090 17900 31100
rect 20940 31260 21100 31270
rect 20940 31090 21100 31100
rect 10620 30480 10700 30490
rect 10620 30370 10700 30380
rect 13320 30480 13420 30490
rect 16080 30480 16180 30490
rect 16080 30370 16180 30380
rect 18820 30480 18920 30490
rect 13320 30350 13420 30360
rect 18820 30350 18920 30360
rect 10580 27920 10760 29040
rect 11660 28780 11820 28790
rect 11660 28310 11820 28320
rect 13300 28140 13460 29040
rect 14360 28780 14520 28790
rect 14360 28310 14520 28320
rect 16060 28140 16220 29040
rect 16480 28780 16640 28790
rect 16480 28310 16640 28320
rect 17120 28780 17280 28790
rect 17120 28310 17280 28320
rect 13300 28020 14440 28140
rect 10580 27820 14040 27920
rect 13880 27620 14040 27820
rect 14280 27620 14440 28020
rect 14700 28020 16220 28140
rect 14700 27620 14840 28020
rect 18800 27920 18960 29040
rect 19860 28780 20020 28790
rect 19860 28310 20020 28320
rect 15080 27820 18960 27920
rect 15080 27620 15240 27820
rect 22740 25860 23740 26020
rect 23600 24080 23740 25860
rect 18440 24020 18580 24030
rect 15040 23980 17880 24000
rect 15040 23860 17520 23980
rect 17620 23860 17880 23980
rect 23600 23940 23880 24080
rect 18440 23870 18580 23880
rect 15040 23840 17880 23860
rect 24940 23680 25080 23690
rect 23260 23660 24020 23680
rect 23260 23580 23280 23660
rect 23360 23580 24020 23660
rect 23260 23560 24020 23580
rect 24940 23550 25080 23560
rect 13420 23380 13540 23390
rect 13420 22230 13540 22240
rect 23500 23160 23880 23320
rect 9320 21780 9680 21790
rect 23500 21740 23680 23160
rect 9320 21610 9680 21620
rect 21300 21560 23680 21740
rect 17740 21380 17860 21390
rect 17740 21250 17860 21260
rect 18760 21360 18860 21370
rect 18760 21250 18860 21260
rect 16020 20220 17940 20230
rect 16020 20050 17940 20060
<< via2 >>
rect 14560 43740 14640 43820
rect 15680 43480 15760 43560
rect 28180 42620 28280 42720
rect 28740 42100 28840 42200
rect 14560 36920 14640 37000
rect 15560 34900 15640 34980
rect 9540 31100 9680 31400
rect 12240 31100 12400 31400
rect 15000 31100 15160 31400
rect 17740 31100 17900 31400
rect 20940 31100 21100 31260
rect 10620 30380 10700 30480
rect 13320 30360 13420 30480
rect 16080 30380 16180 30480
rect 18820 30360 18920 30480
rect 11660 28320 11820 28780
rect 14360 28320 14520 28780
rect 16480 28320 16640 28780
rect 17120 28320 17280 28780
rect 19860 28320 20020 28780
rect 17520 23860 17620 23980
rect 18440 23880 18580 24020
rect 23280 23580 23360 23660
rect 24940 23560 25080 23680
rect 13420 22240 13540 23380
rect 9320 21620 9680 21780
rect 17740 21260 17860 21380
rect 18760 21260 18860 21360
rect 16020 20060 17940 20220
<< metal3 >>
rect 13620 44100 13740 44120
rect 13620 44020 13640 44100
rect 13720 44020 13740 44100
rect 13620 38800 13740 44020
rect 14540 43820 14780 43840
rect 14540 43740 14560 43820
rect 14640 43740 14680 43820
rect 14760 43740 14780 43820
rect 14540 43720 14780 43740
rect 15660 43560 15900 43580
rect 15660 43480 15680 43560
rect 15760 43480 15800 43560
rect 15880 43480 15900 43560
rect 15660 43460 15900 43480
rect 17640 42780 17760 42800
rect 17640 42700 17660 42780
rect 17740 42700 17760 42780
rect 17640 40620 17760 42700
rect 28170 42720 28290 42725
rect 28170 42620 28180 42720
rect 28280 42620 28290 42720
rect 28170 42615 28290 42620
rect 28730 42200 28850 42205
rect 28730 42100 28740 42200
rect 28840 42100 28850 42200
rect 28730 42095 28850 42100
rect 10600 38680 17080 38800
rect 9530 31400 9690 31405
rect 9530 31100 9540 31400
rect 9680 31100 9690 31400
rect 9530 31095 9690 31100
rect 10600 30480 10720 38680
rect 14540 37000 14660 37020
rect 14540 36920 14560 37000
rect 14640 36920 14660 37000
rect 14540 36900 14660 36920
rect 13300 36780 17120 36900
rect 12230 31400 12410 31405
rect 12230 31100 12240 31400
rect 12400 31100 12410 31400
rect 12230 31095 12410 31100
rect 10600 30380 10620 30480
rect 10700 30380 10720 30480
rect 10600 30340 10720 30380
rect 13300 30480 13440 36780
rect 25040 36760 25420 36920
rect 15540 34980 17120 35000
rect 15540 34900 15560 34980
rect 15640 34900 17120 34980
rect 15540 34880 17120 34900
rect 14990 31400 15170 31405
rect 14990 31100 15000 31400
rect 15160 31100 15170 31400
rect 14990 31095 15170 31100
rect 13300 30360 13320 30480
rect 13420 30360 13440 30480
rect 16060 30480 16200 34880
rect 17070 33000 17080 33080
rect 17160 33000 17170 33080
rect 17520 32580 17700 33100
rect 17520 32480 18920 32580
rect 18800 31600 18920 32480
rect 18800 31500 23380 31600
rect 17730 31400 17910 31405
rect 17730 31100 17740 31400
rect 17900 31100 17910 31400
rect 17730 31095 17910 31100
rect 16060 30380 16080 30480
rect 16180 30380 16200 30480
rect 16060 30360 16200 30380
rect 18800 30480 18940 31500
rect 20930 31260 21110 31265
rect 20930 31100 20940 31260
rect 21100 31100 21110 31260
rect 20930 31095 21110 31100
rect 18800 30360 18820 30480
rect 18920 30360 18940 30480
rect 13300 30340 13440 30360
rect 18800 30340 18940 30360
rect 280 28800 9180 28820
rect 280 28300 300 28800
rect 580 28780 22798 28800
rect 580 28320 11660 28780
rect 11820 28320 14360 28780
rect 14520 28320 16480 28780
rect 16640 28320 17120 28780
rect 17280 28320 19860 28780
rect 20020 28770 22798 28780
rect 20020 28327 22005 28770
rect 22334 28327 22798 28770
rect 20020 28320 22798 28327
rect 580 28300 22798 28320
rect 280 28280 9160 28300
rect 9300 21780 9700 28300
rect 18420 24020 21880 24040
rect 17500 23980 17640 24000
rect 17500 23860 17520 23980
rect 17620 23860 17640 23980
rect 18420 23880 18440 24020
rect 18580 23880 21880 24020
rect 18420 23860 21880 23880
rect 13410 23380 13550 23385
rect 13410 22240 13420 23380
rect 13540 22240 13550 23380
rect 13410 22235 13550 22240
rect 9300 21620 9320 21780
rect 9680 21620 9700 21780
rect 9300 21600 9700 21620
rect 17500 21400 17640 23860
rect 17500 21380 17880 21400
rect 17500 21260 17740 21380
rect 17860 21260 17880 21380
rect 17500 21240 17880 21260
rect 18740 21360 18880 21380
rect 18740 21260 18760 21360
rect 18860 21260 18880 21360
rect 16010 20220 17950 20225
rect 16010 20060 16020 20220
rect 17940 20060 17950 20220
rect 16010 20055 17950 20060
rect 18740 18840 18880 21260
rect 21740 18840 21880 23860
rect 23260 23660 23380 31500
rect 25260 23700 25420 36760
rect 23260 23580 23280 23660
rect 23360 23580 23380 23660
rect 23260 23560 23380 23580
rect 24920 23680 25420 23700
rect 24920 23560 24940 23680
rect 25080 23560 25420 23680
rect 24920 23540 25420 23560
rect 18740 18820 30540 18840
rect 18740 18660 30380 18820
rect 30520 18660 30540 18820
rect 18740 18640 30540 18660
<< via3 >>
rect 13640 44020 13720 44100
rect 14680 43740 14760 43820
rect 15800 43480 15880 43560
rect 17660 42700 17740 42780
rect 28180 42620 28280 42720
rect 28740 42100 28840 42200
rect 9540 31100 9680 31400
rect 12240 31100 12400 31400
rect 15000 31100 15160 31400
rect 17080 33000 17160 33080
rect 17740 31100 17900 31400
rect 20940 31100 21100 31260
rect 300 28300 580 28800
rect 22005 28327 22334 28770
rect 13420 22240 13540 23380
rect 16020 20060 17940 20220
rect 30380 18660 30520 18820
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44980 16682 45152
rect 17174 44980 17234 45152
rect 17726 44980 17786 45152
rect 200 28800 600 44152
rect 200 28300 300 28800
rect 580 28300 600 28800
rect 200 1000 600 28300
rect 800 31420 1200 44152
rect 16600 44120 16700 44980
rect 13620 44100 16700 44120
rect 13620 44020 13640 44100
rect 13720 44020 16700 44100
rect 13620 44000 16700 44020
rect 17160 43840 17240 44980
rect 14660 43820 17240 43840
rect 14660 43740 14680 43820
rect 14760 43740 17240 43820
rect 14660 43720 17240 43740
rect 17720 43580 17800 44980
rect 18278 44960 18338 45152
rect 18830 44960 18890 45152
rect 15780 43560 17800 43580
rect 15780 43480 15800 43560
rect 15880 43480 17800 43560
rect 15780 43460 17800 43480
rect 18260 43180 18360 44960
rect 16620 43060 18360 43180
rect 16620 33100 16720 43060
rect 17640 42780 17800 42800
rect 18820 42780 18900 44960
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44980 28274 45152
rect 28766 44980 28826 45152
rect 17640 42700 17660 42780
rect 17740 42700 18900 42780
rect 28200 42740 28280 44980
rect 17640 42680 18900 42700
rect 28160 42720 28300 42740
rect 28160 42620 28180 42720
rect 28280 42620 28300 42720
rect 28160 42600 28300 42620
rect 28740 42220 28840 44980
rect 29318 44952 29378 45152
rect 28720 42200 28860 42220
rect 28720 42100 28740 42200
rect 28840 42100 28860 42200
rect 28720 42080 28860 42100
rect 16620 33080 17180 33100
rect 16620 33000 17080 33080
rect 17160 33000 17180 33080
rect 16620 32980 17180 33000
rect 800 31400 17960 31420
rect 800 31100 9540 31400
rect 9680 31100 12240 31400
rect 12400 31100 15000 31400
rect 15160 31100 17740 31400
rect 17900 31280 17960 31400
rect 19711 31280 20108 34012
rect 17900 31260 21140 31280
rect 17900 31100 20940 31260
rect 21100 31100 21140 31260
rect 800 31080 21140 31100
rect 800 20240 1200 31080
rect 21972 28770 22365 34014
rect 21972 28327 22005 28770
rect 22334 28327 22365 28770
rect 21972 28300 22365 28327
rect 13380 23380 13560 23400
rect 13380 22240 13420 23380
rect 13540 22240 13560 23380
rect 13380 20240 13560 22240
rect 800 20220 18020 20240
rect 800 20060 16020 20220
rect 17940 20060 18020 20220
rect 800 20040 18020 20060
rect 800 1000 1200 20040
rect 30355 18820 30553 18857
rect 30355 18660 30380 18820
rect 30520 18660 30553 18820
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30355 185 30553 18660
rect 30362 0 30542 185
use ART  ART_0
timestamp 1740063090
transform 1 0 4814 0 1 8228
box -2000 -6200 14900 1200
use Comp_Sel  Comp_Sel_0
timestamp 1739975917
transform 1 0 22845 0 1 24511
box 1012 -2269 2266 506
use DAC  DAC_0
timestamp 1739900237
transform 1 0 14685 0 -1 25577
box -1445 -2206 620 3537
use DAC_driver  DAC_driver_0
timestamp 1739891334
transform 0 1 10675 -1 0 31449
box 759 -1182 2458 1185
use DAC_driver  DAC_driver_1
timestamp 1739891334
transform 0 1 13381 -1 0 31444
box 759 -1182 2458 1185
use DAC_driver  DAC_driver_2
timestamp 1739891334
transform 0 1 16142 -1 0 31444
box 759 -1182 2458 1185
use DAC_driver  DAC_driver_3
timestamp 1739891334
transform 0 1 18880 -1 0 31444
box 759 -1182 2458 1185
use NComp  NComp_0
timestamp 1739911419
transform 1 0 16224 0 1 23280
box -299 -3281 5084 -118
use PComp  PComp_0
timestamp 1739974557
transform 1 0 14662 0 -1 26038
box 2398 -1502 8203 2241
use SAR  SAR_0
timestamp 1740303368
transform 1 0 17066 0 1 31880
box 0 0 8127 10271
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
